GENERATOR
Time=0 reset=0  counter=0 count=0 
DRIVER
Time=0 reset=0  counter=0 count=0 
MONITOR
Time=5 reset=0  counter=0 count=0 
SCOREBOARD
Time=5 reset=0  counter=0 count=0 
---------COUNTER IS RESETED--------------
GENERATOR
Time=5 reset=0  counter=1 count=0 
DRIVER
Time=5 reset=0  counter=1 count=0 
MONITOR
Time=15 reset=1  counter=1 count=1 
SCOREBOARD
Time=15 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=15 reset=0  counter=0 count=0 
DRIVER
Time=15 reset=0  counter=0 count=0 
MONITOR
Time=25 reset=1  counter=0 count=0 
SCOREBOARD
Time=25 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=25 reset=0  counter=0 count=0 
DRIVER
Time=25 reset=0  counter=0 count=0 
MONITOR
Time=35 reset=1  counter=0 count=127 
SCOREBOARD
Time=35 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=35 reset=0  counter=1 count=0 
DRIVER
Time=35 reset=0  counter=1 count=0 
MONITOR
Time=45 reset=1  counter=1 count=0 
SCOREBOARD
Time=45 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=45 reset=0  counter=1 count=0 
DRIVER
Time=45 reset=0  counter=1 count=0 
MONITOR
Time=55 reset=1  counter=1 count=1 
SCOREBOARD
Time=55 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=55 reset=0  counter=1 count=0 
DRIVER
Time=55 reset=0  counter=1 count=0 
MONITOR
Time=65 reset=1  counter=1 count=2 
SCOREBOARD
Time=65 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=65 reset=0  counter=1 count=0 
DRIVER
Time=65 reset=0  counter=1 count=0 
MONITOR
Time=75 reset=1  counter=1 count=3 
SCOREBOARD
Time=75 reset=1  counter=1 count=3 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=75 reset=0  counter=0 count=0 
DRIVER
Time=75 reset=0  counter=0 count=0 
MONITOR
Time=85 reset=1  counter=0 count=2 
SCOREBOARD
Time=85 reset=1  counter=0 count=2 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=85 reset=0  counter=1 count=0 
DRIVER
Time=85 reset=0  counter=1 count=0 
MONITOR
Time=95 reset=1  counter=1 count=3 
SCOREBOARD
Time=95 reset=1  counter=1 count=3 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=95 reset=0  counter=0 count=0 
DRIVER
Time=95 reset=0  counter=0 count=0 
MONITOR
Time=105 reset=1  counter=0 count=2 
SCOREBOARD
Time=105 reset=1  counter=0 count=2 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=105 reset=0  counter=0 count=0 
DRIVER
Time=105 reset=0  counter=0 count=0 
MONITOR
Time=115 reset=1  counter=0 count=1 
SCOREBOARD
Time=115 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=115 reset=0  counter=1 count=0 
DRIVER
Time=115 reset=0  counter=1 count=0 
MONITOR
Time=125 reset=1  counter=1 count=2 
SCOREBOARD
Time=125 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=125 reset=0  counter=0 count=0 
DRIVER
Time=125 reset=0  counter=0 count=0 
MONITOR
Time=135 reset=1  counter=0 count=1 
SCOREBOARD
Time=135 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=135 reset=0  counter=0 count=0 
DRIVER
Time=135 reset=0  counter=0 count=0 
MONITOR
Time=145 reset=1  counter=0 count=0 
SCOREBOARD
Time=145 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=145 reset=0  counter=1 count=0 
DRIVER
Time=145 reset=0  counter=1 count=0 
MONITOR
Time=155 reset=1  counter=1 count=1 
SCOREBOARD
Time=155 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=155 reset=0  counter=0 count=0 
DRIVER
Time=155 reset=0  counter=0 count=0 
MONITOR
Time=165 reset=1  counter=0 count=0 
SCOREBOARD
Time=165 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=165 reset=0  counter=1 count=0 
DRIVER
Time=165 reset=0  counter=1 count=0 
MONITOR
Time=175 reset=1  counter=1 count=1 
SCOREBOARD
Time=175 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=175 reset=0  counter=0 count=0 
DRIVER
Time=175 reset=0  counter=0 count=0 
MONITOR
Time=185 reset=1  counter=0 count=0 
SCOREBOARD
Time=185 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=185 reset=0  counter=1 count=0 
DRIVER
Time=185 reset=0  counter=1 count=0 
MONITOR
Time=195 reset=1  counter=1 count=1 
SCOREBOARD
Time=195 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=195 reset=0  counter=1 count=0 
DRIVER
Time=195 reset=0  counter=1 count=0 
MONITOR
Time=205 reset=1  counter=1 count=2 
SCOREBOARD
Time=205 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=205 reset=0  counter=0 count=0 
DRIVER
Time=205 reset=0  counter=0 count=0 
MONITOR
Time=215 reset=1  counter=0 count=1 
SCOREBOARD
Time=215 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=215 reset=0  counter=0 count=0 
DRIVER
Time=215 reset=0  counter=0 count=0 
MONITOR
Time=225 reset=1  counter=0 count=0 
SCOREBOARD
Time=225 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=225 reset=0  counter=0 count=0 
DRIVER
Time=225 reset=0  counter=0 count=0 
MONITOR
Time=235 reset=1  counter=0 count=127 
SCOREBOARD
Time=235 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=235 reset=0  counter=0 count=0 
DRIVER
Time=235 reset=0  counter=0 count=0 
MONITOR
Time=245 reset=1  counter=0 count=126 
SCOREBOARD
Time=245 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=245 reset=0  counter=0 count=0 
DRIVER
Time=245 reset=0  counter=0 count=0 
MONITOR
Time=255 reset=1  counter=0 count=125 
SCOREBOARD
Time=255 reset=1  counter=0 count=125 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=255 reset=0  counter=1 count=0 
DRIVER
Time=255 reset=0  counter=1 count=0 
MONITOR
Time=265 reset=1  counter=1 count=126 
SCOREBOARD
Time=265 reset=1  counter=1 count=126 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=265 reset=0  counter=1 count=0 
DRIVER
Time=265 reset=0  counter=1 count=0 
MONITOR
Time=275 reset=1  counter=1 count=127 
SCOREBOARD
Time=275 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=275 reset=0  counter=1 count=0 
DRIVER
Time=275 reset=0  counter=1 count=0 
MONITOR
Time=285 reset=1  counter=1 count=0 
SCOREBOARD
Time=285 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=285 reset=0  counter=1 count=0 
DRIVER
Time=285 reset=0  counter=1 count=0 
MONITOR
Time=295 reset=1  counter=1 count=1 
SCOREBOARD
Time=295 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=295 reset=0  counter=0 count=0 
DRIVER
Time=295 reset=0  counter=0 count=0 
MONITOR
Time=305 reset=1  counter=0 count=0 
SCOREBOARD
Time=305 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=305 reset=0  counter=0 count=0 
DRIVER
Time=305 reset=0  counter=0 count=0 
MONITOR
Time=315 reset=1  counter=0 count=127 
SCOREBOARD
Time=315 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=315 reset=0  counter=0 count=0 
DRIVER
Time=315 reset=0  counter=0 count=0 
MONITOR
Time=325 reset=1  counter=0 count=126 
SCOREBOARD
Time=325 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=325 reset=0  counter=1 count=0 
DRIVER
Time=325 reset=0  counter=1 count=0 
MONITOR
Time=335 reset=1  counter=1 count=127 
SCOREBOARD
Time=335 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=335 reset=0  counter=0 count=0 
DRIVER
Time=335 reset=0  counter=0 count=0 
MONITOR
Time=345 reset=1  counter=0 count=126 
SCOREBOARD
Time=345 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=345 reset=0  counter=0 count=0 
DRIVER
Time=345 reset=0  counter=0 count=0 
MONITOR
Time=355 reset=1  counter=0 count=125 
SCOREBOARD
Time=355 reset=1  counter=0 count=125 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=355 reset=0  counter=1 count=0 
DRIVER
Time=355 reset=0  counter=1 count=0 
MONITOR
Time=365 reset=1  counter=1 count=126 
SCOREBOARD
Time=365 reset=1  counter=1 count=126 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=365 reset=0  counter=0 count=0 
DRIVER
Time=365 reset=0  counter=0 count=0 
MONITOR
Time=375 reset=1  counter=0 count=125 
SCOREBOARD
Time=375 reset=1  counter=0 count=125 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=375 reset=0  counter=1 count=0 
DRIVER
Time=375 reset=0  counter=1 count=0 
MONITOR
Time=385 reset=1  counter=1 count=126 
SCOREBOARD
Time=385 reset=1  counter=1 count=126 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=385 reset=0  counter=1 count=0 
DRIVER
Time=385 reset=0  counter=1 count=0 
MONITOR
Time=395 reset=1  counter=1 count=127 
SCOREBOARD
Time=395 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=395 reset=0  counter=1 count=0 
DRIVER
Time=395 reset=0  counter=1 count=0 
MONITOR
Time=405 reset=1  counter=1 count=0 
SCOREBOARD
Time=405 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=405 reset=0  counter=0 count=0 
DRIVER
Time=405 reset=0  counter=0 count=0 
MONITOR
Time=415 reset=1  counter=0 count=127 
SCOREBOARD
Time=415 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=415 reset=0  counter=0 count=0 
DRIVER
Time=415 reset=0  counter=0 count=0 
MONITOR
Time=425 reset=1  counter=0 count=126 
SCOREBOARD
Time=425 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=425 reset=0  counter=1 count=0 
DRIVER
Time=425 reset=0  counter=1 count=0 
MONITOR
Time=435 reset=1  counter=1 count=127 
SCOREBOARD
Time=435 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=435 reset=0  counter=0 count=0 
DRIVER
Time=435 reset=0  counter=0 count=0 
MONITOR
Time=445 reset=1  counter=0 count=126 
SCOREBOARD
Time=445 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=445 reset=0  counter=1 count=0 
DRIVER
Time=445 reset=0  counter=1 count=0 
MONITOR
Time=455 reset=1  counter=1 count=127 
SCOREBOARD
Time=455 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=455 reset=0  counter=1 count=0 
DRIVER
Time=455 reset=0  counter=1 count=0 
MONITOR
Time=465 reset=1  counter=1 count=0 
SCOREBOARD
Time=465 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=465 reset=0  counter=0 count=0 
DRIVER
Time=465 reset=0  counter=0 count=0 
MONITOR
Time=475 reset=1  counter=0 count=127 
SCOREBOARD
Time=475 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=475 reset=0  counter=0 count=0 
DRIVER
Time=475 reset=0  counter=0 count=0 
MONITOR
Time=485 reset=1  counter=0 count=126 
SCOREBOARD
Time=485 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=485 reset=0  counter=1 count=0 
DRIVER
Time=485 reset=0  counter=1 count=0 
MONITOR
Time=495 reset=1  counter=1 count=127 
SCOREBOARD
Time=495 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=495 reset=0  counter=1 count=0 
DRIVER
Time=495 reset=0  counter=1 count=0 
MONITOR
Time=505 reset=1  counter=1 count=0 
SCOREBOARD
Time=505 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=505 reset=0  counter=1 count=0 
DRIVER
Time=505 reset=0  counter=1 count=0 
MONITOR
Time=515 reset=1  counter=1 count=1 
SCOREBOARD
Time=515 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=515 reset=0  counter=1 count=0 
DRIVER
Time=515 reset=0  counter=1 count=0 
MONITOR
Time=525 reset=1  counter=1 count=2 
SCOREBOARD
Time=525 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=525 reset=0  counter=0 count=0 
DRIVER
Time=525 reset=0  counter=0 count=0 
MONITOR
Time=535 reset=1  counter=0 count=1 
SCOREBOARD
Time=535 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=535 reset=0  counter=0 count=0 
DRIVER
Time=535 reset=0  counter=0 count=0 
MONITOR
Time=545 reset=1  counter=0 count=0 
SCOREBOARD
Time=545 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=545 reset=0  counter=1 count=0 
DRIVER
Time=545 reset=0  counter=1 count=0 
MONITOR
Time=555 reset=1  counter=1 count=1 
SCOREBOARD
Time=555 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=555 reset=0  counter=1 count=0 
DRIVER
Time=555 reset=0  counter=1 count=0 
MONITOR
Time=565 reset=1  counter=1 count=2 
SCOREBOARD
Time=565 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=565 reset=0  counter=0 count=0 
DRIVER
Time=565 reset=0  counter=0 count=0 
MONITOR
Time=575 reset=1  counter=0 count=1 
SCOREBOARD
Time=575 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=575 reset=0  counter=1 count=0 
DRIVER
Time=575 reset=0  counter=1 count=0 
MONITOR
Time=585 reset=1  counter=1 count=2 
SCOREBOARD
Time=585 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=585 reset=0  counter=0 count=0 
DRIVER
Time=585 reset=0  counter=0 count=0 
MONITOR
Time=595 reset=1  counter=0 count=1 
SCOREBOARD
Time=595 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=595 reset=0  counter=1 count=0 
DRIVER
Time=595 reset=0  counter=1 count=0 
MONITOR
Time=605 reset=1  counter=1 count=2 
SCOREBOARD
Time=605 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=605 reset=0  counter=0 count=0 
DRIVER
Time=605 reset=0  counter=0 count=0 
MONITOR
Time=615 reset=1  counter=0 count=1 
SCOREBOARD
Time=615 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=615 reset=0  counter=0 count=0 
DRIVER
Time=615 reset=0  counter=0 count=0 
MONITOR
Time=625 reset=1  counter=0 count=0 
SCOREBOARD
Time=625 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=625 reset=0  counter=1 count=0 
DRIVER
Time=625 reset=0  counter=1 count=0 
MONITOR
Time=635 reset=1  counter=1 count=1 
SCOREBOARD
Time=635 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=635 reset=0  counter=0 count=0 
DRIVER
Time=635 reset=0  counter=0 count=0 
MONITOR
Time=645 reset=1  counter=0 count=0 
SCOREBOARD
Time=645 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=645 reset=0  counter=1 count=0 
DRIVER
Time=645 reset=0  counter=1 count=0 
MONITOR
Time=655 reset=1  counter=1 count=1 
SCOREBOARD
Time=655 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=655 reset=0  counter=1 count=0 
DRIVER
Time=655 reset=0  counter=1 count=0 
MONITOR
Time=665 reset=1  counter=1 count=2 
SCOREBOARD
Time=665 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=665 reset=0  counter=0 count=0 
DRIVER
Time=665 reset=0  counter=0 count=0 
MONITOR
Time=675 reset=1  counter=0 count=1 
SCOREBOARD
Time=675 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=675 reset=0  counter=0 count=0 
DRIVER
Time=675 reset=0  counter=0 count=0 
MONITOR
Time=685 reset=1  counter=0 count=0 
SCOREBOARD
Time=685 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=685 reset=0  counter=1 count=0 
DRIVER
Time=685 reset=0  counter=1 count=0 
MONITOR
Time=695 reset=1  counter=1 count=1 
SCOREBOARD
Time=695 reset=1  counter=1 count=1 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=695 reset=0  counter=1 count=0 
DRIVER
Time=695 reset=0  counter=1 count=0 
MONITOR
Time=705 reset=1  counter=1 count=2 
SCOREBOARD
Time=705 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=705 reset=0  counter=0 count=0 
DRIVER
Time=705 reset=0  counter=0 count=0 
MONITOR
Time=715 reset=1  counter=0 count=1 
SCOREBOARD
Time=715 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=715 reset=0  counter=1 count=0 
DRIVER
Time=715 reset=0  counter=1 count=0 
MONITOR
Time=725 reset=1  counter=1 count=2 
SCOREBOARD
Time=725 reset=1  counter=1 count=2 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=725 reset=0  counter=1 count=0 
DRIVER
Time=725 reset=0  counter=1 count=0 
MONITOR
Time=735 reset=1  counter=1 count=3 
SCOREBOARD
Time=735 reset=1  counter=1 count=3 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=735 reset=0  counter=1 count=0 
DRIVER
Time=735 reset=0  counter=1 count=0 
MONITOR
Time=745 reset=1  counter=1 count=4 
SCOREBOARD
Time=745 reset=1  counter=1 count=4 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=745 reset=0  counter=0 count=0 
DRIVER
Time=745 reset=0  counter=0 count=0 
MONITOR
Time=755 reset=1  counter=0 count=3 
SCOREBOARD
Time=755 reset=1  counter=0 count=3 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=755 reset=0  counter=0 count=0 
DRIVER
Time=755 reset=0  counter=0 count=0 
MONITOR
Time=765 reset=1  counter=0 count=2 
SCOREBOARD
Time=765 reset=1  counter=0 count=2 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=765 reset=0  counter=1 count=0 
DRIVER
Time=765 reset=0  counter=1 count=0 
MONITOR
Time=775 reset=1  counter=1 count=3 
SCOREBOARD
Time=775 reset=1  counter=1 count=3 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=775 reset=0  counter=0 count=0 
DRIVER
Time=775 reset=0  counter=0 count=0 
MONITOR
Time=785 reset=1  counter=0 count=2 
SCOREBOARD
Time=785 reset=1  counter=0 count=2 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=785 reset=0  counter=0 count=0 
DRIVER
Time=785 reset=0  counter=0 count=0 
MONITOR
Time=795 reset=1  counter=0 count=1 
SCOREBOARD
Time=795 reset=1  counter=0 count=1 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=795 reset=0  counter=0 count=0 
DRIVER
Time=795 reset=0  counter=0 count=0 
MONITOR
Time=805 reset=1  counter=0 count=0 
SCOREBOARD
Time=805 reset=1  counter=0 count=0 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=805 reset=0  counter=0 count=0 
DRIVER
Time=805 reset=0  counter=0 count=0 
MONITOR
Time=815 reset=1  counter=0 count=127 
SCOREBOARD
Time=815 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=815 reset=0  counter=1 count=0 
DRIVER
Time=815 reset=0  counter=1 count=0 
MONITOR
Time=825 reset=1  counter=1 count=0 
SCOREBOARD
Time=825 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=825 reset=0  counter=0 count=0 
DRIVER
Time=825 reset=0  counter=0 count=0 
MONITOR
Time=835 reset=1  counter=0 count=127 
SCOREBOARD
Time=835 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=835 reset=0  counter=0 count=0 
DRIVER
Time=835 reset=0  counter=0 count=0 
MONITOR
Time=845 reset=1  counter=0 count=126 
SCOREBOARD
Time=845 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=845 reset=0  counter=1 count=0 
DRIVER
Time=845 reset=0  counter=1 count=0 
MONITOR
Time=855 reset=1  counter=1 count=127 
SCOREBOARD
Time=855 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=855 reset=0  counter=1 count=0 
DRIVER
Time=855 reset=0  counter=1 count=0 
MONITOR
Time=865 reset=1  counter=1 count=0 
SCOREBOARD
Time=865 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=865 reset=0  counter=0 count=0 
DRIVER
Time=865 reset=0  counter=0 count=0 
MONITOR
Time=875 reset=1  counter=0 count=127 
SCOREBOARD
Time=875 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=875 reset=0  counter=1 count=0 
DRIVER
Time=875 reset=0  counter=1 count=0 
MONITOR
Time=885 reset=1  counter=1 count=0 
SCOREBOARD
Time=885 reset=1  counter=1 count=0 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=885 reset=0  counter=0 count=0 
DRIVER
Time=885 reset=0  counter=0 count=0 
MONITOR
Time=895 reset=1  counter=0 count=127 
SCOREBOARD
Time=895 reset=1  counter=0 count=127 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=895 reset=0  counter=0 count=0 
DRIVER
Time=895 reset=0  counter=0 count=0 
MONITOR
Time=905 reset=1  counter=0 count=126 
SCOREBOARD
Time=905 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=905 reset=0  counter=1 count=0 
DRIVER
Time=905 reset=0  counter=1 count=0 
MONITOR
Time=915 reset=1  counter=1 count=127 
SCOREBOARD
Time=915 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=915 reset=0  counter=0 count=0 
DRIVER
Time=915 reset=0  counter=0 count=0 
MONITOR
Time=925 reset=1  counter=0 count=126 
SCOREBOARD
Time=925 reset=1  counter=0 count=126 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=925 reset=0  counter=0 count=0 
DRIVER
Time=925 reset=0  counter=0 count=0 
MONITOR
Time=935 reset=1  counter=0 count=125 
SCOREBOARD
Time=935 reset=1  counter=0 count=125 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=935 reset=0  counter=0 count=0 
DRIVER
Time=935 reset=0  counter=0 count=0 
MONITOR
Time=945 reset=1  counter=0 count=124 
SCOREBOARD
Time=945 reset=1  counter=0 count=124 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=945 reset=0  counter=1 count=0 
DRIVER
Time=945 reset=0  counter=1 count=0 
MONITOR
Time=955 reset=1  counter=1 count=125 
SCOREBOARD
Time=955 reset=1  counter=1 count=125 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=955 reset=0  counter=1 count=0 
DRIVER
Time=955 reset=0  counter=1 count=0 
MONITOR
Time=965 reset=1  counter=1 count=126 
SCOREBOARD
Time=965 reset=1  counter=1 count=126 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=965 reset=0  counter=0 count=0 
DRIVER
Time=965 reset=0  counter=0 count=0 
MONITOR
Time=975 reset=1  counter=0 count=125 
SCOREBOARD
Time=975 reset=1  counter=0 count=125 
----------DOWNCOUNTER IS PASSED-------------- 
GENERATOR
Time=975 reset=0  counter=1 count=0 
DRIVER
Time=975 reset=0  counter=1 count=0 
MONITOR
Time=985 reset=1  counter=1 count=126 
SCOREBOARD
Time=985 reset=1  counter=1 count=126 
----------UPCOUNTER IS PASSED-------------- 
GENERATOR
Time=985 reset=0  counter=1 count=0 
DRIVER
Time=985 reset=0  counter=1 count=0 
MONITOR
Time=995 reset=1  counter=1 count=127 
SCOREBOARD
Time=995 reset=1  counter=1 count=127 
----------UPCOUNTER IS PASSED-------------- 
$finish at simulation time                  995
