GENERATOR
data_in=1000 sel=1 data_out=0 
DRIVER
data_in=1000 sel=1 data_out=0 
MONITOR
data_in=1000 sel=1 data_out=1100 
SCOREBOARD
data_in=1000 sel=1 data_out=1100 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=1001 sel=1 data_out=0 
DRIVER
data_in=1001 sel=1 data_out=0 
MONITOR
data_in=1001 sel=1 data_out=1101 
SCOREBOARD
data_in=1001 sel=1 data_out=1101 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=0 sel=1 data_out=0 
DRIVER
data_in=0 sel=1 data_out=0 
MONITOR
data_in=0 sel=1 data_out=0 
SCOREBOARD
data_in=0 sel=1 data_out=0 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=1000 sel=1 data_out=0 
DRIVER
data_in=1000 sel=1 data_out=0 
MONITOR
data_in=1000 sel=1 data_out=1100 
SCOREBOARD
data_in=1000 sel=1 data_out=1100 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=101 sel=1 data_out=0 
DRIVER
data_in=101 sel=1 data_out=0 
MONITOR
data_in=101 sel=1 data_out=111 
SCOREBOARD
data_in=101 sel=1 data_out=111 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=11 sel=1 data_out=0 
DRIVER
data_in=11 sel=1 data_out=0 
MONITOR
data_in=11 sel=1 data_out=10 
SCOREBOARD
data_in=11 sel=1 data_out=10 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=1001 sel=1 data_out=0 
DRIVER
data_in=1001 sel=1 data_out=0 
MONITOR
data_in=1001 sel=1 data_out=1101 
SCOREBOARD
data_in=1001 sel=1 data_out=1101 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=11 sel=1 data_out=0 
DRIVER
data_in=11 sel=1 data_out=0 
MONITOR
data_in=11 sel=1 data_out=10 
SCOREBOARD
data_in=11 sel=1 data_out=10 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=1100 sel=1 data_out=0 
DRIVER
data_in=1100 sel=1 data_out=0 
MONITOR
data_in=1100 sel=1 data_out=1010 
SCOREBOARD
data_in=1100 sel=1 data_out=1010 
PASS----------------binary to gray------------------PASS
GENERATOR
data_in=101 sel=1 data_out=0 
DRIVER
data_in=101 sel=1 data_out=0 
MONITOR
data_in=101 sel=1 data_out=111 
SCOREBOARD
data_in=101 sel=1 data_out=111 
PASS----------------binary to gray------------------PASS
$finish at simulation time                   30
