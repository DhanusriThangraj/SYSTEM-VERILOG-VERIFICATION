interface inter;
  logic [3:0]a;
  logic [3:0]b;
  logic [1:0]sel;
  logic [5:0]sum;
  logic [5:0]sub;
  logic [8:0]mul;
  logic [3:0]div;
endinterface
