GENERATOR
Time=0 reset=0 d=0 q=0
DRIVER
Time=5 reset=0 d=0 q=0
reset=1
MONITOR
Time=5 reset=1 d=0 q=0
SCOREBOARD
Time=5 reset=1 d=0 q=0
---------PASS---------
GENERATOR
Time=5 reset=0 d=1 q=0
MONITOR
Time=15 reset=1 d=0 q=0
DRIVER
Time=15 reset=0 d=1 q=0
reset=1
SCOREBOARD
Time=15 reset=1 d=0 q=0
---------PASS---------
GENERATOR
Time=15 reset=0 d=0 q=0
MONITOR
Time=25 reset=0 d=1 q=1
DRIVER
Time=25 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=25 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=25 reset=0 d=0 q=0
MONITOR
Time=35 reset=0 d=0 q=0
DRIVER
Time=35 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=35 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=35 reset=0 d=1 q=0
MONITOR
Time=45 reset=0 d=0 q=0
DRIVER
Time=45 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=45 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=45 reset=0 d=1 q=0
MONITOR
Time=55 reset=0 d=1 q=1
DRIVER
Time=55 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=55 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=55 reset=0 d=1 q=0
MONITOR
Time=65 reset=0 d=1 q=1
DRIVER
Time=65 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=65 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=65 reset=0 d=1 q=0
MONITOR
Time=75 reset=0 d=1 q=1
DRIVER
Time=75 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=75 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=75 reset=0 d=0 q=0
MONITOR
Time=85 reset=0 d=1 q=1
DRIVER
Time=85 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=85 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=85 reset=0 d=1 q=0
MONITOR
Time=95 reset=0 d=0 q=0
DRIVER
Time=95 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=95 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=95 reset=0 d=0 q=0
MONITOR
Time=105 reset=0 d=1 q=1
DRIVER
Time=105 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=105 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=105 reset=0 d=0 q=0
MONITOR
Time=115 reset=0 d=0 q=0
DRIVER
Time=115 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=115 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=115 reset=0 d=1 q=0
MONITOR
Time=125 reset=0 d=0 q=0
DRIVER
Time=125 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=125 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=125 reset=0 d=0 q=0
MONITOR
Time=135 reset=0 d=1 q=1
DRIVER
Time=135 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=135 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=135 reset=0 d=0 q=0
MONITOR
Time=145 reset=0 d=0 q=0
DRIVER
Time=145 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=145 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=145 reset=0 d=1 q=0
MONITOR
Time=155 reset=0 d=0 q=0
DRIVER
Time=155 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=155 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=155 reset=0 d=0 q=0
MONITOR
Time=165 reset=0 d=1 q=1
DRIVER
Time=165 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=165 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=165 reset=0 d=1 q=0
MONITOR
Time=175 reset=0 d=0 q=0
DRIVER
Time=175 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=175 reset=0 d=0 q=0
---------PASS---------
GENERATOR
Time=175 reset=0 d=0 q=0
MONITOR
Time=185 reset=0 d=1 q=1
DRIVER
Time=185 reset=0 d=0 q=0
reset=0
SCOREBOARD
Time=185 reset=0 d=1 q=1
---------PASS---------
GENERATOR
Time=185 reset=0 d=1 q=0
MONITOR
Time=195 reset=0 d=0 q=0
DRIVER
Time=195 reset=0 d=1 q=0
reset=0
SCOREBOARD
Time=195 reset=0 d=0 q=0
---------PASS---------
