interface inter;
  logic [3:0]data_in;
  logic sel;
  logic [3:0]data_out;
endinterface
