GENERATOR
 Time=0 a=0 b=1 c=1 sum=0 carry=0
DRIVER
 Time=1 a=0 b=1 c=1 sum=0 carry=0
MONITOR
 Time=2 a=0 b=1 c=1 sum=0 carry=1
SCOREBOARD
 Time=2 a=0 b=1 c=1 sum=0 carry=1
===================PASS======================
SCOREBOARD
 Time=2 a=0 b=1 c=1 sum=0 carry=1
GENERATOR
 Time=3 a=1 b=1 c=1 sum=0 carry=0
DRIVER
 Time=4 a=1 b=1 c=1 sum=0 carry=0
MONITOR
 Time=5 a=1 b=1 c=1 sum=1 carry=1
SCOREBOARD
 Time=5 a=1 b=1 c=1 sum=1 carry=1
===================PASS======================
SCOREBOARD
 Time=5 a=1 b=1 c=1 sum=1 carry=1
$finish at simulation time     
