GENERATOR
TIME=0 reset=0 din=9 addr=15 en=1 dout=0
DRIVER
TIME=0 reset=0 din=9 addr=15 en=1 dout=0
MONITOR
TIME=5 reset=1 din=9 addr=15 en=1 dout=0
SCOREBOARD
TIME=5 reset=1 din=9 addr=15 en=1 dout=0
----------------RAM MEMORY IS RESETED----------------
GENERATOR
TIME=5 reset=0 din=13 addr=11 en=1 dout=0
DRIVER
TIME=5 reset=0 din=13 addr=11 en=1 dout=0
MONITOR
TIME=15 reset=1 din=13 addr=11 en=1 dout=0
SCOREBOARD
TIME=15 reset=1 din=13 addr=11 en=1 dout=0
----------------RAM MEMORY IS RESETED----------------
GENERATOR
TIME=15 reset=0 din=9 addr=0 en=1 dout=0
DRIVER
TIME=15 reset=0 din=9 addr=0 en=1 dout=0
MONITOR
TIME=25 reset=1 din=9 addr=0 en=1 dout=0
SCOREBOARD
TIME=25 reset=1 din=9 addr=0 en=1 dout=0
----------------RAM MEMORY IS RESETED----------------
GENERATOR
TIME=25 reset=0 din=1 addr=13 en=0 dout=0
DRIVER
TIME=25 reset=0 din=1 addr=13 en=0 dout=0
MONITOR
TIME=35 reset=1 din=1 addr=13 en=0 dout=0
SCOREBOARD
TIME=35 reset=1 din=1 addr=13 en=0 dout=0
----------------RAM MEMORY IS RESETED----------------
GENERATOR
TIME=35 reset=0 din=10 addr=6 en=1 dout=0
DRIVER
TIME=35 reset=0 din=10 addr=6 en=1 dout=0
MONITOR
TIME=45 reset=0 din=10 addr=6 en=1 dout=0
SCOREBOARD
TIME=45 reset=0 din=10 addr=6 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=45 reset=0 din=1 addr=11 en=0 dout=0
DRIVER
TIME=45 reset=0 din=1 addr=11 en=0 dout=0
MONITOR
TIME=55 reset=0 din=1 addr=11 en=0 dout=0
SCOREBOARD
TIME=55 reset=0 din=1 addr=11 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=55 reset=0 din=9 addr=2 en=1 dout=0
DRIVER
TIME=55 reset=0 din=9 addr=2 en=1 dout=0
MONITOR
TIME=65 reset=0 din=9 addr=2 en=1 dout=0
SCOREBOARD
TIME=65 reset=0 din=9 addr=2 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=65 reset=0 din=3 addr=3 en=0 dout=0
DRIVER
TIME=65 reset=0 din=3 addr=3 en=0 dout=0
MONITOR
TIME=75 reset=0 din=3 addr=3 en=0 dout=0
SCOREBOARD
TIME=75 reset=0 din=3 addr=3 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=75 reset=0 din=11 addr=9 en=1 dout=0
DRIVER
TIME=75 reset=0 din=11 addr=9 en=1 dout=0
MONITOR
TIME=85 reset=0 din=11 addr=9 en=1 dout=0
SCOREBOARD
TIME=85 reset=0 din=11 addr=9 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=85 reset=0 din=3 addr=3 en=0 dout=0
DRIVER
TIME=85 reset=0 din=3 addr=3 en=0 dout=0
MONITOR
TIME=95 reset=0 din=3 addr=3 en=0 dout=0
SCOREBOARD
TIME=95 reset=0 din=3 addr=3 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=95 reset=0 din=15 addr=10 en=0 dout=0
DRIVER
TIME=95 reset=0 din=15 addr=10 en=0 dout=0
MONITOR
TIME=105 reset=0 din=15 addr=10 en=0 dout=0
SCOREBOARD
TIME=105 reset=0 din=15 addr=10 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=105 reset=0 din=5 addr=15 en=1 dout=0
DRIVER
TIME=105 reset=0 din=5 addr=15 en=1 dout=0
MONITOR
TIME=115 reset=0 din=5 addr=15 en=1 dout=0
SCOREBOARD
TIME=115 reset=0 din=5 addr=15 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=115 reset=0 din=5 addr=11 en=0 dout=0
DRIVER
TIME=115 reset=0 din=5 addr=11 en=0 dout=0
MONITOR
TIME=125 reset=0 din=5 addr=11 en=0 dout=0
SCOREBOARD
TIME=125 reset=0 din=5 addr=11 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=125 reset=0 din=9 addr=0 en=0 dout=0
DRIVER
TIME=125 reset=0 din=9 addr=0 en=0 dout=0
MONITOR
TIME=135 reset=0 din=9 addr=0 en=0 dout=0
SCOREBOARD
TIME=135 reset=0 din=9 addr=0 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=135 reset=0 din=3 addr=7 en=0 dout=0
DRIVER
TIME=135 reset=0 din=3 addr=7 en=0 dout=0
MONITOR
TIME=145 reset=0 din=3 addr=7 en=0 dout=0
SCOREBOARD
TIME=145 reset=0 din=3 addr=7 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=145 reset=0 din=8 addr=1 en=1 dout=0
DRIVER
TIME=145 reset=0 din=8 addr=1 en=1 dout=0
MONITOR
TIME=155 reset=0 din=8 addr=1 en=1 dout=0
SCOREBOARD
TIME=155 reset=0 din=8 addr=1 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=155 reset=0 din=13 addr=1 en=0 dout=0
DRIVER
TIME=155 reset=0 din=13 addr=1 en=0 dout=0
MONITOR
TIME=165 reset=0 din=13 addr=1 en=0 dout=8
SCOREBOARD
TIME=165 reset=0 din=13 addr=1 en=0 dout=8
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=165 reset=0 din=14 addr=1 en=0 dout=0
DRIVER
TIME=165 reset=0 din=14 addr=1 en=0 dout=0
MONITOR
TIME=175 reset=0 din=14 addr=1 en=0 dout=8
SCOREBOARD
TIME=175 reset=0 din=14 addr=1 en=0 dout=8
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=175 reset=0 din=14 addr=1 en=0 dout=0
DRIVER
TIME=175 reset=0 din=14 addr=1 en=0 dout=0
MONITOR
TIME=185 reset=0 din=14 addr=1 en=0 dout=8
SCOREBOARD
TIME=185 reset=0 din=14 addr=1 en=0 dout=8
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=185 reset=0 din=14 addr=1 en=0 dout=0
DRIVER
TIME=185 reset=0 din=14 addr=1 en=0 dout=0
MONITOR
TIME=195 reset=0 din=14 addr=1 en=0 dout=8
SCOREBOARD
TIME=195 reset=0 din=14 addr=1 en=0 dout=8
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=195 reset=0 din=5 addr=11 en=0 dout=0
DRIVER
TIME=195 reset=0 din=5 addr=11 en=0 dout=0
MONITOR
TIME=205 reset=0 din=5 addr=11 en=0 dout=0
SCOREBOARD
TIME=205 reset=0 din=5 addr=11 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=205 reset=0 din=14 addr=5 en=0 dout=0
DRIVER
TIME=205 reset=0 din=14 addr=5 en=0 dout=0
MONITOR
TIME=215 reset=0 din=14 addr=5 en=0 dout=0
SCOREBOARD
TIME=215 reset=0 din=14 addr=5 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=215 reset=0 din=6 addr=10 en=1 dout=0
DRIVER
TIME=215 reset=0 din=6 addr=10 en=1 dout=0
MONITOR
TIME=225 reset=0 din=6 addr=10 en=1 dout=0
SCOREBOARD
TIME=225 reset=0 din=6 addr=10 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=225 reset=0 din=9 addr=0 en=0 dout=0
DRIVER
TIME=225 reset=0 din=9 addr=0 en=0 dout=0
MONITOR
TIME=235 reset=0 din=9 addr=0 en=0 dout=0
SCOREBOARD
TIME=235 reset=0 din=9 addr=0 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=235 reset=0 din=8 addr=0 en=1 dout=0
DRIVER
TIME=235 reset=0 din=8 addr=0 en=1 dout=0
MONITOR
TIME=245 reset=0 din=8 addr=0 en=1 dout=0
SCOREBOARD
TIME=245 reset=0 din=8 addr=0 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=245 reset=0 din=13 addr=7 en=1 dout=0
DRIVER
TIME=245 reset=0 din=13 addr=7 en=1 dout=0
MONITOR
TIME=255 reset=0 din=13 addr=7 en=1 dout=0
SCOREBOARD
TIME=255 reset=0 din=13 addr=7 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=255 reset=0 din=0 addr=15 en=1 dout=0
DRIVER
TIME=255 reset=0 din=0 addr=15 en=1 dout=0
MONITOR
TIME=265 reset=0 din=0 addr=15 en=1 dout=0
SCOREBOARD
TIME=265 reset=0 din=0 addr=15 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=265 reset=0 din=11 addr=15 en=0 dout=0
DRIVER
TIME=265 reset=0 din=11 addr=15 en=0 dout=0
MONITOR
TIME=275 reset=0 din=11 addr=15 en=0 dout=0
SCOREBOARD
TIME=275 reset=0 din=11 addr=15 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=275 reset=0 din=13 addr=13 en=1 dout=0
DRIVER
TIME=275 reset=0 din=13 addr=13 en=1 dout=0
MONITOR
TIME=285 reset=0 din=13 addr=13 en=1 dout=0
SCOREBOARD
TIME=285 reset=0 din=13 addr=13 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=285 reset=0 din=10 addr=5 en=1 dout=0
DRIVER
TIME=285 reset=0 din=10 addr=5 en=1 dout=0
MONITOR
TIME=295 reset=0 din=10 addr=5 en=1 dout=0
SCOREBOARD
TIME=295 reset=0 din=10 addr=5 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=295 reset=0 din=8 addr=8 en=0 dout=0
DRIVER
TIME=295 reset=0 din=8 addr=8 en=0 dout=0
MONITOR
TIME=305 reset=0 din=8 addr=8 en=0 dout=0
SCOREBOARD
TIME=305 reset=0 din=8 addr=8 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=305 reset=0 din=12 addr=11 en=1 dout=0
DRIVER
TIME=305 reset=0 din=12 addr=11 en=1 dout=0
MONITOR
TIME=315 reset=0 din=12 addr=11 en=1 dout=0
SCOREBOARD
TIME=315 reset=0 din=12 addr=11 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=315 reset=0 din=4 addr=8 en=0 dout=0
DRIVER
TIME=315 reset=0 din=4 addr=8 en=0 dout=0
MONITOR
TIME=325 reset=0 din=4 addr=8 en=0 dout=0
SCOREBOARD
TIME=325 reset=0 din=4 addr=8 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=325 reset=0 din=6 addr=2 en=1 dout=0
DRIVER
TIME=325 reset=0 din=6 addr=2 en=1 dout=0
MONITOR
TIME=335 reset=0 din=6 addr=2 en=1 dout=0
SCOREBOARD
TIME=335 reset=0 din=6 addr=2 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=335 reset=0 din=8 addr=0 en=0 dout=0
DRIVER
TIME=335 reset=0 din=8 addr=0 en=0 dout=0
MONITOR
TIME=345 reset=0 din=8 addr=0 en=0 dout=8
SCOREBOARD
TIME=345 reset=0 din=8 addr=0 en=0 dout=8
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=345 reset=0 din=13 addr=14 en=0 dout=0
DRIVER
TIME=345 reset=0 din=13 addr=14 en=0 dout=0
MONITOR
TIME=355 reset=0 din=13 addr=14 en=0 dout=0
SCOREBOARD
TIME=355 reset=0 din=13 addr=14 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=355 reset=0 din=3 addr=12 en=1 dout=0
DRIVER
TIME=355 reset=0 din=3 addr=12 en=1 dout=0
MONITOR
TIME=365 reset=0 din=3 addr=12 en=1 dout=0
SCOREBOARD
TIME=365 reset=0 din=3 addr=12 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=365 reset=0 din=2 addr=3 en=1 dout=0
DRIVER
TIME=365 reset=0 din=2 addr=3 en=1 dout=0
MONITOR
TIME=375 reset=0 din=2 addr=3 en=1 dout=0
SCOREBOARD
TIME=375 reset=0 din=2 addr=3 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=375 reset=0 din=3 addr=12 en=0 dout=0
DRIVER
TIME=375 reset=0 din=3 addr=12 en=0 dout=0
MONITOR
TIME=385 reset=0 din=3 addr=12 en=0 dout=3
SCOREBOARD
TIME=385 reset=0 din=3 addr=12 en=0 dout=3
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=385 reset=0 din=11 addr=2 en=1 dout=0
DRIVER
TIME=385 reset=0 din=11 addr=2 en=1 dout=0
MONITOR
TIME=395 reset=0 din=11 addr=2 en=1 dout=3
SCOREBOARD
TIME=395 reset=0 din=11 addr=2 en=1 dout=3
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=395 reset=0 din=0 addr=0 en=1 dout=0
DRIVER
TIME=395 reset=0 din=0 addr=0 en=1 dout=0
MONITOR
TIME=405 reset=0 din=0 addr=0 en=1 dout=3
SCOREBOARD
TIME=405 reset=0 din=0 addr=0 en=1 dout=3
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=405 reset=0 din=11 addr=15 en=0 dout=0
DRIVER
TIME=405 reset=0 din=11 addr=15 en=0 dout=0
MONITOR
TIME=415 reset=0 din=11 addr=15 en=0 dout=0
SCOREBOARD
TIME=415 reset=0 din=11 addr=15 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=415 reset=0 din=13 addr=2 en=1 dout=0
DRIVER
TIME=415 reset=0 din=13 addr=2 en=1 dout=0
MONITOR
TIME=425 reset=0 din=13 addr=2 en=1 dout=0
SCOREBOARD
TIME=425 reset=0 din=13 addr=2 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=425 reset=0 din=2 addr=15 en=1 dout=0
DRIVER
TIME=425 reset=0 din=2 addr=15 en=1 dout=0
MONITOR
TIME=435 reset=0 din=2 addr=15 en=1 dout=0
SCOREBOARD
TIME=435 reset=0 din=2 addr=15 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=435 reset=0 din=6 addr=5 en=0 dout=0
DRIVER
TIME=435 reset=0 din=6 addr=5 en=0 dout=0
MONITOR
TIME=445 reset=0 din=6 addr=5 en=0 dout=10
SCOREBOARD
TIME=445 reset=0 din=6 addr=5 en=0 dout=10
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=445 reset=0 din=12 addr=15 en=1 dout=0
DRIVER
TIME=445 reset=0 din=12 addr=15 en=1 dout=0
MONITOR
TIME=455 reset=0 din=12 addr=15 en=1 dout=10
SCOREBOARD
TIME=455 reset=0 din=12 addr=15 en=1 dout=10
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=455 reset=0 din=8 addr=9 en=1 dout=0
DRIVER
TIME=455 reset=0 din=8 addr=9 en=1 dout=0
MONITOR
TIME=465 reset=0 din=8 addr=9 en=1 dout=10
SCOREBOARD
TIME=465 reset=0 din=8 addr=9 en=1 dout=10
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=465 reset=0 din=3 addr=2 en=0 dout=0
DRIVER
TIME=465 reset=0 din=3 addr=2 en=0 dout=0
MONITOR
TIME=475 reset=0 din=3 addr=2 en=0 dout=13
SCOREBOARD
TIME=475 reset=0 din=3 addr=2 en=0 dout=13
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=475 reset=0 din=15 addr=9 en=1 dout=0
DRIVER
TIME=475 reset=0 din=15 addr=9 en=1 dout=0
MONITOR
TIME=485 reset=0 din=15 addr=9 en=1 dout=13
SCOREBOARD
TIME=485 reset=0 din=15 addr=9 en=1 dout=13
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=485 reset=0 din=1 addr=15 en=0 dout=0
DRIVER
TIME=485 reset=0 din=1 addr=15 en=0 dout=0
MONITOR
TIME=495 reset=0 din=1 addr=15 en=0 dout=12
SCOREBOARD
TIME=495 reset=0 din=1 addr=15 en=0 dout=12
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=495 reset=0 din=13 addr=1 en=1 dout=0
DRIVER
TIME=495 reset=0 din=13 addr=1 en=1 dout=0
MONITOR
TIME=505 reset=0 din=13 addr=1 en=1 dout=12
SCOREBOARD
TIME=505 reset=0 din=13 addr=1 en=1 dout=12
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=505 reset=0 din=10 addr=9 en=1 dout=0
DRIVER
TIME=505 reset=0 din=10 addr=9 en=1 dout=0
MONITOR
TIME=515 reset=0 din=10 addr=9 en=1 dout=12
SCOREBOARD
TIME=515 reset=0 din=10 addr=9 en=1 dout=12
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=515 reset=0 din=5 addr=11 en=1 dout=0
DRIVER
TIME=515 reset=0 din=5 addr=11 en=1 dout=0
MONITOR
TIME=525 reset=0 din=5 addr=11 en=1 dout=12
SCOREBOARD
TIME=525 reset=0 din=5 addr=11 en=1 dout=12
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=525 reset=0 din=0 addr=8 en=0 dout=0
DRIVER
TIME=525 reset=0 din=0 addr=8 en=0 dout=0
MONITOR
TIME=535 reset=0 din=0 addr=8 en=0 dout=0
SCOREBOARD
TIME=535 reset=0 din=0 addr=8 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=535 reset=0 din=7 addr=9 en=1 dout=0
DRIVER
TIME=535 reset=0 din=7 addr=9 en=1 dout=0
MONITOR
TIME=545 reset=0 din=7 addr=9 en=1 dout=0
SCOREBOARD
TIME=545 reset=0 din=7 addr=9 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=545 reset=0 din=0 addr=7 en=1 dout=0
DRIVER
TIME=545 reset=0 din=0 addr=7 en=1 dout=0
MONITOR
TIME=555 reset=0 din=0 addr=7 en=1 dout=0
SCOREBOARD
TIME=555 reset=0 din=0 addr=7 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=555 reset=0 din=14 addr=14 en=0 dout=0
DRIVER
TIME=555 reset=0 din=14 addr=14 en=0 dout=0
MONITOR
TIME=565 reset=0 din=14 addr=14 en=0 dout=0
SCOREBOARD
TIME=565 reset=0 din=14 addr=14 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=565 reset=0 din=3 addr=7 en=1 dout=0
DRIVER
TIME=565 reset=0 din=3 addr=7 en=1 dout=0
MONITOR
TIME=575 reset=0 din=3 addr=7 en=1 dout=0
SCOREBOARD
TIME=575 reset=0 din=3 addr=7 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=575 reset=0 din=5 addr=7 en=1 dout=0
DRIVER
TIME=575 reset=0 din=5 addr=7 en=1 dout=0
MONITOR
TIME=585 reset=0 din=5 addr=7 en=1 dout=0
SCOREBOARD
TIME=585 reset=0 din=5 addr=7 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=585 reset=0 din=6 addr=5 en=0 dout=0
DRIVER
TIME=585 reset=0 din=6 addr=5 en=0 dout=0
MONITOR
TIME=595 reset=0 din=6 addr=5 en=0 dout=10
SCOREBOARD
TIME=595 reset=0 din=6 addr=5 en=0 dout=10
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=595 reset=0 din=11 addr=9 en=1 dout=0
DRIVER
TIME=595 reset=0 din=11 addr=9 en=1 dout=0
MONITOR
TIME=605 reset=0 din=11 addr=9 en=1 dout=10
SCOREBOARD
TIME=605 reset=0 din=11 addr=9 en=1 dout=10
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=605 reset=0 din=15 addr=6 en=1 dout=0
DRIVER
TIME=605 reset=0 din=15 addr=6 en=1 dout=0
MONITOR
TIME=615 reset=0 din=15 addr=6 en=1 dout=10
SCOREBOARD
TIME=615 reset=0 din=15 addr=6 en=1 dout=10
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=615 reset=0 din=15 addr=1 en=0 dout=0
DRIVER
TIME=615 reset=0 din=15 addr=1 en=0 dout=0
MONITOR
TIME=625 reset=0 din=15 addr=1 en=0 dout=13
SCOREBOARD
TIME=625 reset=0 din=15 addr=1 en=0 dout=13
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=625 reset=0 din=11 addr=8 en=0 dout=0
DRIVER
TIME=625 reset=0 din=11 addr=8 en=0 dout=0
MONITOR
TIME=635 reset=0 din=11 addr=8 en=0 dout=0
SCOREBOARD
TIME=635 reset=0 din=11 addr=8 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=635 reset=0 din=0 addr=6 en=0 dout=0
DRIVER
TIME=635 reset=0 din=0 addr=6 en=0 dout=0
MONITOR
TIME=645 reset=0 din=0 addr=6 en=0 dout=15
SCOREBOARD
TIME=645 reset=0 din=0 addr=6 en=0 dout=15
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=645 reset=0 din=15 addr=9 en=1 dout=0
DRIVER
TIME=645 reset=0 din=15 addr=9 en=1 dout=0
MONITOR
TIME=655 reset=0 din=15 addr=9 en=1 dout=15
SCOREBOARD
TIME=655 reset=0 din=15 addr=9 en=1 dout=15
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=655 reset=0 din=13 addr=15 en=0 dout=0
DRIVER
TIME=655 reset=0 din=13 addr=15 en=0 dout=0
MONITOR
TIME=665 reset=0 din=13 addr=15 en=0 dout=12
SCOREBOARD
TIME=665 reset=0 din=13 addr=15 en=0 dout=12
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=665 reset=0 din=8 addr=9 en=1 dout=0
DRIVER
TIME=665 reset=0 din=8 addr=9 en=1 dout=0
MONITOR
TIME=675 reset=0 din=8 addr=9 en=1 dout=12
SCOREBOARD
TIME=675 reset=0 din=8 addr=9 en=1 dout=12
----------------DATA WRITE IS PASSED----------------
GENERATOR
TIME=675 reset=0 din=13 addr=8 en=0 dout=0
DRIVER
TIME=675 reset=0 din=13 addr=8 en=0 dout=0
MONITOR
TIME=685 reset=0 din=13 addr=8 en=0 dout=0
SCOREBOARD
TIME=685 reset=0 din=13 addr=8 en=0 dout=0
----------------DATA READ IS PASSED----------------
GENERATOR
TIME=685 reset=0 din=7 addr=7 en=1 dout=0
DRIVER
TIME=685 reset=0 din=7 addr=7 en=1 dout=0
MONITOR
TIME=695 reset=0 din=7 addr=7 en=1 dout=0
SCOREBOARD
TIME=695 reset=0 din=7 addr=7 en=1 dout=0
----------------DATA WRITE IS PASSED----------------
