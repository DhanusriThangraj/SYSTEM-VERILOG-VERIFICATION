GENERATOR
Time=0 a=8 b=9 sel=3 sum=0 sub=0 mul=0 div=0
DRIVER
Time=1 a=8 b=9 sel=3 sum=0 sub=0 mul=0 div=0
MONITOR
Time=2 a=8 b=9 sel=3 sum=0 sub=0 mul=0 div=0
SCOREBOARD
Time=2 a=8 b=9 sel=3 sum=0 sub=0 mul=0 div=0
DIV-----------PASS------------DIV
GENERATOR
Time=3 a=9 b=3 sel=1 sum=0 sub=0 mul=0 div=0
DRIVER
Time=4 a=9 b=3 sel=1 sum=0 sub=0 mul=0 div=0
MONITOR
Time=5 a=9 b=3 sel=1 sum=0 sub=6 mul=0 div=0
SCOREBOARD
Time=5 a=9 b=3 sel=1 sum=0 sub=6 mul=0 div=0
SUB-----------PASS------------SUB
GENERATOR
Time=6 a=0 b=3 sel=3 sum=0 sub=0 mul=0 div=0
DRIVER
Time=7 a=0 b=3 sel=3 sum=0 sub=0 mul=0 div=0
MONITOR
Time=8 a=0 b=3 sel=3 sum=0 sub=6 mul=0 div=0
SCOREBOARD
Time=8 a=0 b=3 sel=3 sum=0 sub=6 mul=0 div=0
DIV-----------PASS------------DIV
GENERATOR
Time=9 a=8 b=13 sel=0 sum=0 sub=0 mul=0 div=0
DRIVER
Time=10 a=8 b=13 sel=0 sum=0 sub=0 mul=0 div=0
MONITOR
Time=11 a=8 b=13 sel=0 sum=21 sub=6 mul=0 div=0
SCOREBOARD
Time=11 a=8 b=13 sel=0 sum=21 sub=6 mul=0 div=0
SUM-----------PASS------------SUM
GENERATOR
Time=12 a=5 b=11 sel=0 sum=0 sub=0 mul=0 div=0
DRIVER
Time=13 a=5 b=11 sel=0 sum=0 sub=0 mul=0 div=0
MONITOR
Time=14 a=5 b=11 sel=0 sum=16 sub=6 mul=0 div=0
SCOREBOARD
Time=14 a=5 b=11 sel=0 sum=16 sub=6 mul=0 div=0
SUM-----------PASS------------SUM
GENERATOR
Time=15 a=3 b=7 sel=2 sum=0 sub=0 mul=0 div=0
DRIVER
Time=16 a=3 b=7 sel=2 sum=0 sub=0 mul=0 div=0
MONITOR
Time=17 a=3 b=7 sel=2 sum=16 sub=6 mul=21 div=0
SCOREBOARD
Time=17 a=3 b=7 sel=2 sum=16 sub=6 mul=21 div=0
MUL-----------PASS------------MUL
GENERATOR
Time=18 a=9 b=13 sel=3 sum=0 sub=0 mul=0 div=0
DRIVER
Time=19 a=9 b=13 sel=3 sum=0 sub=0 mul=0 div=0
MONITOR
Time=20 a=9 b=13 sel=3 sum=16 sub=6 mul=21 div=0
SCOREBOARD
Time=20 a=9 b=13 sel=3 sum=16 sub=6 mul=21 div=0
DIV-----------PASS------------DIV
GENERATOR
Time=21 a=3 b=5 sel=1 sum=0 sub=0 mul=0 div=0
DRIVER
Time=22 a=3 b=5 sel=1 sum=0 sub=0 mul=0 div=0
MONITOR
Time=23 a=3 b=5 sel=1 sum=16 sub=-2 mul=21 div=0
SCOREBOARD
Time=23 a=3 b=5 sel=1 sum=16 sub=-2 mul=21 div=0
SUB-----------PASS------------SUB
GENERATOR
Time=24 a=12 b=1 sel=0 sum=0 sub=0 mul=0 div=0
DRIVER
Time=25 a=12 b=1 sel=0 sum=0 sub=0 mul=0 div=0
MONITOR
Time=26 a=12 b=1 sel=0 sum=13 sub=-2 mul=21 div=0
SCOREBOARD
Time=26 a=12 b=1 sel=0 sum=13 sub=-2 mul=21 div=0
SUM-----------PASS------------SUM
GENERATOR
Time=27 a=5 b=15 sel=3 sum=0 sub=0 mul=0 div=0
DRIVER
Time=28 a=5 b=15 sel=3 sum=0 sub=0 mul=0 div=0
MONITOR
Time=29 a=5 b=15 sel=3 sum=13 sub=-2 mul=21 div=0
SCOREBOARD
Time=29 a=5 b=15 sel=3 sum=13 sub=-2 mul=21 div=0
DIV-----------PASS------------DIV
GENERATOR
Time=30 a=14 b=7 sel=1 sum=0 sub=0 mul=0 div=0
DRIVER
Time=31 a=14 b=7 sel=1 sum=0 sub=0 mul=0 div=0
MONITOR
Time=32 a=14 b=7 sel=1 sum=13 sub=7 mul=21 div=0
SCOREBOARD
Time=32 a=14 b=7 sel=1 sum=13 sub=7 mul=21 div=0
SUB-----------PASS------------SUB
GENERATOR
Time=33 a=10 b=2 sel=1 sum=0 sub=0 mul=0 div=0
DRIVER
Time=34 a=10 b=2 sel=1 sum=0 sub=0 mul=0 div=0
MONITOR
Time=35 a=10 b=2 sel=1 sum=13 sub=8 mul=21 div=0
SCOREBOARD
Time=35 a=10 b=2 sel=1 sum=13 sub=8 mul=21 div=0
SUB-----------PASS------------SUB
$finish at simulation time                   
