GENERATOR
Time=0 a=0 b=1 sum=0 carry=0
DRIVER
Time=1 a=0 b=1 sum=0 carry=0
MONITOR
Time=2 a=0 b=1 sum=1 carry=0
SCOREBOARD
Time=2 a=0 b=1 sum=1 carry=0
PASS---------------------------PASS
GENERATOR
Time=3 a=1 b=1 sum=0 carry=0
DRIVER
Time=4 a=1 b=1 sum=0 carry=0
MONITOR
Time=5 a=1 b=1 sum=0 carry=1
SCOREBOARD
Time=5 a=1 b=1 sum=0 carry=1
PASS---------------------------PASS
GENERATOR
Time=6 a=0 b=1 sum=0 carry=0
DRIVER
Time=7 a=0 b=1 sum=0 carry=0
MONITOR
Time=8 a=0 b=1 sum=1 carry=0
SCOREBOARD
Time=8 a=0 b=1 sum=1 carry=0
PASS---------------------------PASS
GENERATOR
Time=9 a=0 b=1 sum=0 carry=0
DRIVER
Time=10 a=0 b=1 sum=0 carry=0
MONITOR
Time=11 a=0 b=1 sum=1 carry=0
SCOREBOARD
Time=11 a=0 b=1 sum=1 carry=0
PASS---------------------------PASS
GENERATOR
Time=12 a=1 b=1 sum=0 carry=0
DRIVER
Time=13 a=1 b=1 sum=0 carry=0
MONITOR
Time=14 a=1 b=1 sum=0 carry=1
SCOREBOARD
Time=14 a=1 b=1 sum=0 carry=1
PASS---------------------------PASS
$finish at simulation time                   15
