interface inter();
  logic clk;
  logic reset;
  logic counter;
  logic [6:0]count;  
endinterface
